`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NUS ECE
// Engineer: Shahzor Ahmad
// 
// Create Date: 02.10.2015 14:31:19
// Design Name: 
// Module Name: SCOPE_TOP
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module SCOPE_TOP(

    input CLK,                  // main system clock, 100MHz
        
    input btnL,                 // buttons
    input btnR,    
    input btnU,
    input btnD,
    
    input ADC_IN_P,             // differential +ve & -ve analog inputs to ADC
    input ADC_IN_N,  
    input triggerSwitch,
    input shiftYSwitch,
    
    output reg[3:0] VGA_RED,    // RGB outputs to VGA connector (4 bits per channel gives 4096 possible colors)
    output reg[3:0] VGA_GREEN,
    output reg[3:0] VGA_BLUE,
    output reg VGA_VS,          // horizontal & vertical sync outputs to VGA connector
    output reg VGA_HS,
     
    output [15:0] led           // debug LEDs    
    
    );   
         
    //-------------------------------------------------------------------------
    
    wire CLK_MAIN = CLK ;   // this is just a renaming (simply a short-circuit, or two names for the same trace/route)           
       
        
    //-------------------------------------------------------------------------
    
    //         INSTANTITATE EXTERNAL MODULES FOR VGA CONTROL
    
    // Note the VGA controller is configured to produce a 1024 x 1280 pixel resolution
    //-------------------------------------------------------------------------
    
    // PIXEL CLOCK GENERATOR 
    wire CLK_VGA ;          // pixel/VGA clock is generated by MMCM/PLL via external VHDL code (108MHz)    
    clk_wiz_0 PIXEL_CLOCK_GENERATOR( 
            CLK_MAIN,   // 100 MHz
            CLK_VGA     // 108 MHz
        ) ;     
    
    
    // VGA SIGNALS (as output by VGA controller (vga_ctrl.vhd))
    wire VGA_horzSync ;
    wire VGA_vertSync ;
    wire VGA_active ;
    wire[11:0] VGA_horzCoord ;
    wire[11:0] VGA_vertCoord ;
        // it is not required but good practice to declare single-bit wires
        // it is required to declare multi-bit wires (bus) before use    
    
    // VGA CONTROLLER    
    vga_ctrl VGA_CONTROLLER(
            CLK_VGA,
            VGA_horzSync,
            VGA_vertSync,
            VGA_active,  
            VGA_horzCoord,  
            VGA_vertCoord  
        ) ; 
        // - VGA_horzCoord changes at a rate of 108 MHz (CLK_VGA) to traverse each pixel in a row, while VGA_vertCoord changes at a rate of ~63.98 KHz to 
        // scan each row one by one and back to the top. These tech details are handled by vga_ctrl.vhd. One only needs to make use of these coordinates 
        // to output whatever they want at desired pixel locations. 
        // 
        // - VGA_active is a binary indicator specifying when VGA_horzCoord, VGA_vertCoord are valid (i.e., within the 1024 x 1280 pixel screen). For technical 
        // reasons the said coordinates do go outside this screen area for a short while and no VGA signal should be output during this time (it will and does
        // mess up the display). 
        //
        // - hence, VGA_active, VGA_horzCoord and VGA_vertCoord may be used in conjunction with each other to generate VGA_RED, VGA_GREEN, VGA_BLUE. The Sync
        // signals should be output to the VGA port as well, and are responsible to generate the raster scan on the screen       


    //-------------------------------------------------------------------------
                                    
    //                      SAMPLING VIA ADC 
    
    // On-chip ADC is clocked at [ inv(inv(CLK_ADC/4)*26) = 961.538 KHZ ], 
    // where CLK_ADC is the clock passed to ADC (in this case CLK_ADC = CLK_MAIN = 100MHz)
    
    // The on-chip ADC is 12-bit. Let's use only the most significant 8 bits to keep things simple
    
    //-------------------------------------------------------------------------
    
    wire [7:0] ADC_SAMPLE ; // the latest value as sampled via ADC
    ADC_sampler SAMPLER( CLK_MAIN, ADC_IN_P, ADC_IN_N, ADC_SAMPLE ) ; // sampling at 961.538 KHZ
        // EITHER line # 105 OR lines # 129-135 should be used at a time

    assign led[15:8] = ADC_SAMPLE ;
        // the sampled 8-bit value reflects on 8 LEDs. Every time ADC_SAMPLE changes 
        // (and that happens at 961.538KHz!), this assignment is triggered again 
    assign led[7:4] = 4'd0 ; // force low (you may use these LEDs for debug/indication purposes if needed) 
    
    //-------------------------------------------------------------------------
                                        
    //                  SIMULATE SAMPLING VIA ADC 
    
    // In the absence of a signal generator (e.g., when working at home), you may use 
    // the following code instead of the above, i.e., COMMENT out line # 105, 
    // UN-COMMENT lines # 129-135
    
    // A square wave at 1Hz is 'synthesized' via a clock-divider module, and serves as our 
    // 'analog' signal to be sampled.
    //-------------------------------------------------------------------------
    
    wire CLK_SYNTH_SQUARE ; 
    clock_divider GEN_CLK_SYNTH_SQUARE( CLK_MAIN, 1'b0, 28'H2FAF080, CLK_SYNTH_SQUARE ) ; 
        // Synthesize a 1Hz waveform given 100MHz clock          

//    always@(posedge CLK_MAIN) // sample the synthesized waveform at 100 MHz
//        begin
//            if( CLK_SYNTH_SQUARE )
//                ADC_SAMPLE <= 255 ;
//            else
//                ADC_SAMPLE <= 0 ;        
//        end   
        
//      reg dirn = 1;
//      always@(posedge CLK_SUBSAMPLE) // sample the synthesized waveform at 100 MHz
//          begin
//              if (dirn) 
//                  ADC_SAMPLE = ADC_SAMPLE + 1 ; 
//              else
//                  ADC_SAMPLE = ADC_SAMPLE - 1 ;
             
//              if (ADC_SAMPLE == 8'b1111_1111 || ADC_SAMPLE==0) 
//                  dirn=~dirn;   
//          end      
 
     reg LED_DEBUG = 0 ;
        // this LED blinks at 0.5 Hz (just for visualization)
        // recall, signals on LHS of assignments in 'always' blocks must be declared as reg before use
        
     always@(posedge CLK_SYNTH_SQUARE)
        begin
            LED_DEBUG <= ~LED_DEBUG ;
        end

     assign led[0] = LED_DEBUG ; 
        
               
    //-----------------------------------------------------------------------------------------
                                    
    //        SELECTING SAMPLING FREQUENCY (ESSENTIALLY, CONFIGURING OSCILLOSCOPE's TIME/DIV)
    
    // this configures the CLK_SUBSAMPLE (fs)
    
    // NOTE: currently CLK_SUBSAMPLE_ID has been hard-coded to 0, and no provision
    // is made to modify it at FPGA run-time
    //------------------------------------------------------------------------------------------
    
    reg [3:0] CLK_SUBSAMPLE_ID = 7 ; 
    assign led[3:1] = CLK_SUBSAMPLE_ID ;  
        // leds[11:9] provide a visual indication of CLK_SUBSAMPLE_ID at all times    
        
    reg [27:0] LOAD_VALUE_SUBSAMPLE ;
        // we generate CLK_SUBSAMPLE from CLK_MAIN 
    reg [16:0] LOAD_SHIFT_CLOCK_SAMPLE_RATE  = 28'd125000 ;
    
    always@(CLK_SUBSAMPLE_ID)
        case(CLK_SUBSAMPLE_ID)
            0:  LOAD_VALUE_SUBSAMPLE <= 28'd500000 ;    // CLK_SUBSAMPLE = 100 Hz       => TIME/DIV = 0.8 sec/div
            1:  LOAD_VALUE_SUBSAMPLE <= 28'd250000 ;    // CLK_SUBSAMPLE = 200 Hz       => TIME/DIV = 0.4 sec/div
            2:  LOAD_VALUE_SUBSAMPLE <= 28'd125000 ;    // CLK_SUBSAMPLE = 400 Hz       => TIME/DIV = 0.2 sec/div 
            3:  LOAD_VALUE_SUBSAMPLE <= 28'd62500 ;     // CLK_SUBSAMPLE = 800 Hz       => TIME/DIV = 0.1 sec/div
            4:  LOAD_VALUE_SUBSAMPLE <= 28'd50000 ;     // CLK_SUBSAMPLE = 1 KHz        => TIME/DIV = 80 ms/div
            5:  LOAD_VALUE_SUBSAMPLE <= 28'd31250 ;     // CLK_SUBSAMPLE = 1600 Hz      => TIME/DIV = 50 ms/div 
            6:  LOAD_VALUE_SUBSAMPLE <= 28'd6250 ;      // CLK_SUBSAMPLE = 8 KHz        => TIME/DIV = 10 ms/div 
            7:  LOAD_VALUE_SUBSAMPLE <= 28'd625 ;       // CLK_SUBSAMPLE = 80 KHz       => TIME/DIV = 1 ms/div      
            8:  LOAD_VALUE_SUBSAMPLE <= 28'd62 ;        // CLK_SUBSAMPLE = 806.451 KHz  => TIME/DIV = 0.0992 ms/div 
            9:  LOAD_VALUE_SUBSAMPLE <= 28'd50 ;        // CLK_SUBSAMPLE = 1 MHz        => TIME/DIV = 0.08 ms/div
            10: LOAD_VALUE_SUBSAMPLE <= 28'd6 ;         // CLK_SUBSAMPLE = 8 MHz        => TIME/DIV = 0.01 ms/div
        endcase
            // notice, this is a simple combinational circuit -- for every possible input combination, there's a defined/hard-coded output
            // Each LOAD_VALUE_SUBSAMPLE defines the stated CLK_SUBSAMPLE (sampling frequency fs). 
            // The TIME/DIV values, however, assume the 1280 horizontal pixels on the screen are divided into 16 equal DIVISIONS of 80 px each 
                        
    wire CLK_SUBSAMPLE ;    // sub-sampling rate for ADC output samples
                            // It essentially defines time/div 
                            
                            // Use CLK_SUBSAMPLE to clock your bank of shift registers below
                            // Use CLK_SUBSAMPLE to clock your triggering process when you implement one   
                            
                            // For all practical purposes, this can be taken to be our fs (sampling frequency) as described in the manual
                            // We could have modified ADC sampling frequency, but given the long formula to dervie it from CLK_MAIN (see line 97),
                            // we're better off fixing it, and instead using a sub-sampling frequency to achieve flexible sampling frequencies 
                            // and corresponding time/div configurations
                                                        
                                                     
    clock_divider GEN_CLK_SUBSAMPLE( CLK_MAIN, 1'b0, LOAD_VALUE_SUBSAMPLE, CLK_SUBSAMPLE ) ;
        // note: as many times you instantiate a module in HDL, that many times it will replicate the actual hardware on the FPGA 
        // so this is the 2nd physical clock_divider circuit in our hardware design    
    clock_divider GEN_CLK_SHIFT( CLK_MAIN, 1'b0, LOAD_SHIFT_CLOCK_SAMPLE_RATE, CLK_FOR_SHIFT ) ;
    
    // un-comment lines # 200 - 218 to use PBs to control CLK_SUBSAMPLE_ID, and hence your oscilloscope's TIME/DIV
    // NOTE: you must write Verilog code for a single pulse generator in single_pulse_generator.v for the following to work
    clock_divider GEN_CLK_IN_SINGLE_PULSE( CLK_MAIN, 1'b0, 28'h4C4640, CLK_IN_SINGLE_PULSE ) ;
//        // For CLK_IN_SINGLE_PULSE = 10Hz (100ms), we need LOAD_VALUE = 0d5,000,000 = 0x4C4640 
//        // this would be a 3rd clock-divider in our hardware   

    wire btnL_SINGLE_PULSE ;
    wire btnR_SINGLE_PULSE ; // recall, declaration not needed for single-bit wires, but good practice
    single_pulse_generator btnL_SPG( CLK_IN_SINGLE_PULSE, btnL, btnL_SINGLE_PULSE ) ;
    single_pulse_generator btnR_SPG( CLK_IN_SINGLE_PULSE, btnR, btnR_SINGLE_PULSE ) ;
    single_pulse_generator btnU_SPG( CLK_IN_SINGLE_PULSE, btnU, btnU_SINGLE_PULSE ) ;
    single_pulse_generator btnD_SPG( CLK_IN_SINGLE_PULSE, btnD, btnD_SINGLE_PULSE ) ;
        // note: a separate single pulse generator needs to be instantiated for each push button under use
        // a single_pulse_generator not only provides a single pulse lasting for 1 clock cycle, 
        // but also debounces the switch, killing 2 birds in 1 stone :)
 
    always@(posedge CLK_IN_SINGLE_PULSE) // don't use CLK_MAIN -- the behaviour will then be different from what we intend. Can you explain why?
        begin
            if( btnL_SINGLE_PULSE && CLK_SUBSAMPLE_ID > 0)
                begin
                CLK_SUBSAMPLE_ID <= CLK_SUBSAMPLE_ID - 1 ;
                end
                
            if( btnR_SINGLE_PULSE && CLK_SUBSAMPLE_ID < 10)
                begin
                CLK_SUBSAMPLE_ID <= CLK_SUBSAMPLE_ID + 1 ;
                end
        end
 
    // =============================================>> 
    // CAUTION: Never un-comment the code herein (unless you intend to examine said error). 
    // Use the above version (lines # 212 - 218) instead    
    //
    // the following results in an error ("mult-driven net") during synthesis! 
    // That is, a single physical net/bus (CLK_SUBSAMPLE_ID) will be driven by multiple sources (btnL_SINGLE_PULSE, btnR_SINGLE_PULSE). 
    // In other words, we're short-circuiting two inputs: btnL_SINGLE_PULSE and btnR_SINGLE_PULSE !
    // This was ok in Lab#4 where the output was being driven by only one input, not so here.
    //  
//    always@(posedge btnL_SINGLE_PULSE)
//        begin
//            CLK_SUBSAMPLE_ID = CLK_SUBSAMPLE_ID - 1 ;
//        end
//    always@(posedge btnR_SINGLE_PULSE)
//        begin
//            CLK_SUBSAMPLE_ID = CLK_SUBSAMPLE_ID + 1 ;
//        end
    // ===============================================<<
    
    //-------------------------------------------------------------------------
                                    
    //               UPDATE DISPLAY_MEM @ CLK_SUBSAMPLE
    
    // DISPLAY_MEM is a bank of 1280 shift registers, each 8-bit wide
    //
    // shift all samples one position to the left in memory, and  
    // store the latest ADC sample in the right/left most position    
    //-------------------------------------------------------------------------

    reg [7:0] DISPLAY_MEM[0:1279] ; 
        // display memory - any waveform whose samples are stored here is displayed on screen by the VGA controller
        
    // TOOD:    implement Verilog here that treats DISPLAY_MEM as a bank of 
    //          1280 shift registers, each 8-bit wide. The latest sample should 
    //          be stored in the right (or left)-most register, while contents of
    //          all the other registers should be shifted to the neighboring register
    //          on the right (respectively, left). 
    //          
    //          This process of bringing in a new sample from the right/left while 
    //          shifting all the other samples should be done in a single clock cycle 
    //          (use CLK_SUBSAMPLE)

    reg [10:0] counter;  
    reg [7:0] TEMP_DISPLAY[0:1279] ;
  
    reg squareWave ;
    
    always @(posedge CLK_SUBSAMPLE)
    begin
         if(DISPLAY_MEM[0] == DISPLAY_MEM[1] && DISPLAY_MEM[1] == DISPLAY_MEM[2] && DISPLAY_MEM[2] == DISPLAY_MEM[3] )
            begin
            squareWave <= 1;
            end 
         else
            begin
            squareWave <= 0;
            end
         TEMP_DISPLAY[0] <= ADC_SAMPLE;
     
         for(counter=1; counter < 1280 ; counter = counter +1)
             begin
             TEMP_DISPLAY[counter] <= TEMP_DISPLAY[counter-1];
             end
        
        if(triggerSwitch)
            begin
                       
            if((squareWave && ADC_SAMPLE > 8'd200) || (!squareWave && ADC_SAMPLE > 8'd200 && ADC_SAMPLE < 8'd205 && ADC_SAMPLE < TEMP_DISPLAY[0]))
                begin
                for(counter=1; counter < 1280 ; counter = counter +1)
                    begin
                    DISPLAY_MEM[counter] <= TEMP_DISPLAY[counter]; 
                    end
                end
            end
        else
            begin
        
            for(counter=0; counter < 1280 ; counter = counter +1)
                begin
                DISPLAY_MEM[counter] <= TEMP_DISPLAY[counter];
                end
            end        
    end
    
    
    //-------------------------------------------------------------------------
                
    //                  DRAWING WAVEFORM ON SCREEN
    
    // waveform is drawn using its samples from display memory
    //-------------------------------------------------------------------------       
   
    reg[10:0] yPos = 640;
    always@(posedge CLK_FOR_SHIFT) // don't use CLK_MAIN -- the behaviour will then be different from what we intend. Can you explain why?
            begin
                if( btnU && triggerSwitch && shiftYSwitch && (yPos<1023))
                    begin
                    yPos<= yPos + 1;
                    end
                    
                if( btnD && triggerSwitch && shiftYSwitch && (yPos>255))
                    begin
                    yPos <= yPos - 1;
                    end
            end
    
    
   
                 
    wire[3:0] VGA_WAVEFORM = 
            ((VGA_horzCoord < 1280) & (VGA_vertCoord == (yPos - DISPLAY_MEM[VGA_horzCoord]))) 
                ? 4'hF : 0 ;     
                  
        
    //-------------------------------------------------------------------------
        
    //                  DRAWING GRID LINES ON SCREEN
    
    // Grid lines are drawn at pixels # 320, 640, 960 along the x-axis, and
    // pixels # 256, 512, 768 along the y-axis
    
    // Note the VGA controller is configured to produce a 1024 x 1280 pixel resolution
    //-------------------------------------------------------------------------
            
    wire CONDITION_FOR_GRID = !(VGA_horzCoord % 80) || !(VGA_vertCoord % 64) || ((VGA_horzCoord >= 638)&&(VGA_horzCoord<=642)&&!(VGA_vertCoord % 8))
                                ||((VGA_vertCoord >= 509)&&(VGA_vertCoord<=513)&&!(VGA_horzCoord%16));
    
    wire[3:0] VGA_RED_GRID = CONDITION_FOR_GRID ? 4'hF : 0 ;
    wire[3:0] VGA_GREEN_GRID = CONDITION_FOR_GRID ? 4'hF : 0 ;
    wire[3:0] VGA_BLUE_GRID = CONDITION_FOR_GRID ? 4'hF : 0 ;
        // if true, a black pixel is put at coordinates (VGA_horzCoord, VGA_vertCoord), 
        // else a cyan background is generated, characteristic of oscilloscopes! 
        
    // TOOD:    Draw grid lines at every 80-th pixel along the horizontal axis, and every 64th pixel
    //          along the vertical axis. This gives us a 16x16 grid on screen. 
    //          
    //          Further draw ticks on the central x and y grid lines spaced 16 and 8 pixels apart in the 
    //          horizontal and vertical directions respectively. This gives us 5 sub-divisions per division 
    //          in the horizontal and 8 sub-divisions per divsion in the vertical direction   
    
        
    wire CONDITION_FOR_TIME; 
    CONDITION_TIME conditionTime(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_TIME);                                                                        
    wire[3:0] VGA_TIME = (CONDITION_FOR_TIME)? 4'hF : 0;
    
    wire CONDITION_FOR_SLASH;
    CONDITION_SLASH conditionSlash(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_SLASH);
    wire [3:0] VGA_SLASH = (CONDITION_FOR_SLASH)? 4'hF : 0;
    
    
    wire CONDITION_FOR_COLON = ((VGA_horzCoord == 234) && ((VGA_vertCoord == 943) || (VGA_vertCoord == 947)));  
    wire [3:0] VGA_COLON = (CONDITION_FOR_COLON)? 4'hF : 0;
    
    
    wire CONDITION_FOR_DIV;
    CONDITION_DIV conditionDiv(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_DIV);
    wire [3:0] VGA_DIV = (CONDITION_FOR_DIV)? 4'hF : 0;
    
    wire CONDITION_FOR_FS_0;
    CONDITION_ZERO_EIGHT conditionfs0(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_0);
    
    wire CONDITION_FOR_FS_1;
    CONDITION_FOR_ZERO_FOUR conditionfs1(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_1);
    
    wire CONDITION_FOR_FS_2;
    CONDITION_ZERO_TWO conditionfs2(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_2);
    
    wire CONDITION_FOR_FS_3;
    CONDITION_ZERO_ONE conditionfs3(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_3);
    
    wire CONDITION_FOR_FS_4;
    CONDITION_EIGHT_ZERO_MS conditionfs4(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_4);
    
    wire CONDITION_FOR_FS_5;
    CONDITION_FIFTY_ZERO_MS conditionfs5(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_5);
    
    wire CONDITION_FOR_FS_6;
    CONDITION_ONE_ZERO_MS conditionfs6(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_6);
    
    wire CONDITION_FOR_FS_7;
    CONDITION_ONE_MS conditionfs7(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_7);
    
    wire CONDITION_FOR_FS_8;
    CONDITION_ZERO_ONE_MS conditionfs8(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_8);
    
    wire CONDITION_FOR_FS_9;
    CONDITION_ZERO_ZERO_EIGHT conditionfs9(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_9);
    
    wire CONDITION_FOR_FS_10;
    CONDITION_ZERO_ZERO_ONE_MS conditionfs10(VGA_horzCoord, VGA_vertCoord, CONDITION_FOR_FS_10);
    reg subsampleID_CONDITION;
    always @(CLK_SUBSAMPLE_ID)
        begin
        case (CLK_SUBSAMPLE_ID)
        0:  subsampleID_CONDITION <= CONDITION_FOR_FS_0;
        1:  subsampleID_CONDITION <= CONDITION_FOR_FS_1;
        2:  subsampleID_CONDITION <= CONDITION_FOR_FS_2;
        3:  subsampleID_CONDITION <= CONDITION_FOR_FS_3;
        4:  subsampleID_CONDITION <= CONDITION_FOR_FS_4;
        5:  subsampleID_CONDITION <= CONDITION_FOR_FS_5;
        6:  subsampleID_CONDITION <= CONDITION_FOR_FS_6;
        7:  subsampleID_CONDITION <= CONDITION_FOR_FS_7;
        8:  subsampleID_CONDITION <= CONDITION_FOR_FS_8;
        9:  subsampleID_CONDITION <= CONDITION_FOR_FS_9;
        10: subsampleID_CONDITION <= CONDITION_FOR_FS_10;
        endcase
        end
    
    wire [3:0] VGA_FS = (subsampleID_CONDITION)? 4'hF : 0;
    
    //-------------------------------------------------------------------------
    
    //              SYNCHRONOUS OUTPUT OF VGA SIGNALS
    
    //-------------------------------------------------------------------------
    
    // COMBINE ALL OUTPUTS ON EACH CHANNEL
    wire[3:0] VGA_RED_CHAN = VGA_RED_GRID ;
    wire[3:0] VGA_GREEN_CHAN = VGA_GREEN_GRID | VGA_WAVEFORM | VGA_FS | VGA_TIME | VGA_SLASH | VGA_DIV | VGA_COLON; 
    wire[3:0] VGA_BLUE_CHAN = VGA_BLUE_GRID ;   

    // CLOCK THEM OUT
    always@(posedge CLK_VGA)
        begin      
        
            VGA_RED <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_RED_CHAN ;  
            VGA_GREEN <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_GREEN_CHAN ; 
            VGA_BLUE <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_BLUE_CHAN ; 
                // VGA_active turns off output to screen if scan lines are outside the active screen area
            
            VGA_HS <= VGA_horzSync ;
            VGA_VS <= VGA_vertSync ;
            
        end

    
endmodule
